module top_module(
  input a,
  input b,
  output out
);
  mod_a ma(a, b, out);
endmodule
